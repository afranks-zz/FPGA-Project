
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.all;

package ROMS is
type Sprite is array (0 to 1023) of std_logic_vector(0 to 11);
constant Floor : Sprite := ("101110010110","101110010110","101110010110","100110000100","101010000101","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","011001010011","101110010110","100110000100","100110000100","101110010110","101110010110","100110000100","011001010011","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","011001010011","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","011001010011","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","100110000100","100110000100","101110010110","101110010110","101010000101","100110000100","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","101110010110","101110010110","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","100110000100","100110000100","101110010110","101010000101","101010000101","011001010011","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","011001010011","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","101010000101","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","101110010110","101110010110","100110000100","101110010110","101110010110","101110010110","101110010110","101010000101","100110000100","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","010000110010","010000110010","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011101100011","011101100011","011001010011","011001010011","011001010011","011001010011","011101100011","011101100011","011001010011","011001010011","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","101110010110","101010000101","101010000101","101110010110","100110000100","101110010110","101110010110","101110010110","101110010110","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","101110010110","100110000100","100110000100","100110000100","101110010110","100110000100","100110000100","100110000100","100110000100","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","011001010011","011001010011","100110000100","101110010110","100110000100","100110000100","100110000100","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","011001010011","101010000101","101010000101","101010000101","101010000101","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","101110010110","100110000100","100110000100","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","011001010011","100110000100","100110000100","100110000100","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","011001010011","101010000101","101010000101","101010000101","101110010110","101110010110","101010000101","101010000101","100110000100","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","100110000100","100110000100","100110000100","101010000101","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101110010110","101110010110","101010000101","101010000101","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","100110000100","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","011001010011","011001010011","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101110010110","101110010110","100110000100","101010000101","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","011001010011","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","011001010011","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101010000101","100110000100","100110000100","100110000100","100110000100","100110000100","101010000101","101010000101","101110010110","101110010110","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","101010000101","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","101110010110","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","100110000100","101110010110","101110010110","101110010110","101110010110","101110010110","101010000101","101010000101","101010000101","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","101110010110","100110000100","101110010110","101110010110","100110000100","100110000100","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011","011001010011");
constant BG : Sprite := ("100110011001","101010101010","100110011001","100110011001","101010101010","101010101010","100110011001","101010101010","100010001000","100010001000","101010101010","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","101010101010","100010001000","100010001000","100010001000","100010001000","100010001000","101110111011","010101010101","100010001000","100110011001","101010101010","100110011001","100110011001","101010101010","101010101010","101010101010","101010101010","100010001000","100010001000","101010101010","101010101010","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","100110011001","101010101010","101010101010","100010001000","100010001000","100010001000","100010001000","100110011001","101010101010","010101010101","010101010101","100110011001","100110011001","011101110111","100010001000","100010001000","100010001000","100010001000","100010001000","011001100110","011001100110","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","010101010101","011001100110","101010101010","101010101010","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","011001100110","011001100110","100010001000","100010001000","100010001000","100010001000","100010001000","100110011001","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","011101110111","100010001000","010101010101","011001100110","100010001000","100010001000","011001100110","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","011001100110","011001100110","010101010101","010101010101","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011101110111","011001100110","011001100110","010101010101","010101010101","100110011001","100110011001","011001100110","011001100110","100010001000","011101110111","100110011001","100110011001","011101110111","011101110111","011101110111","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","101010101010","011001100110","011101110111","010101010101","011001100110","100110011001","100110011001","011001100110","011001100110","100010001000","011101110111","100110011001","100110011001","011101110111","011101110111","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","011101110111","011101110111","011101110111","100010001000","100110011001","011001100110","011001100110","010101010101","011001100110","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","100110011001","011001100110","011001100110","011101110111","011101110111","100010001000","100010001000","011101110111","011101110111","010101010101","010101010101","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","100010001000","100110011001","011001100110","011001100110","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","010101010101","010101010101","100010001000","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","011001100110","011001100110","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011101110111","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","010101010101","011001100110","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","011101110111","011101110111","100010001000","100010001000","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","010101010101","010101010101","100010001000","100110011001","011001100110","011001100110","011101110111","011101110111","011001100110","011101110111","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","010101010101","010101010101","011001100110","011001100110","011101110111","011101110111","011101110111","100010001000","010101010101","010101010101","101110111011","101010101010","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","010101010101","011001100110","010101010101","010001000100","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","011001100110","011001100110","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010001000100","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","011001100110","011001100110","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","110011001100","100110011001","101010101010","101010101010","100110011001","100110011001","101010101010","101010101010","101010101010","101010101010","101010101010","101010101010","101110111011","110111011101","010101010101","010101010101","111111111111","110111011101","101010101010","101010101010","101010101010","101110111011","100110011001","100110011001","101010101010","101010101010","101010101010","101110111011","100110011001","100110011001","101110111011","110111011101","101110111011","100110011001","101010101010","100110011001","100110011001","100110011001","100110011001","100110011001","101010101010","101010101010","101010101010","101010101010","101010101010","110111011101","010101010101","010101010101","110111011101","101010101010","100110011001","101010101010","101010101010","101110111011","100110011001","100110011001","101010101010","101010101010","101010101010","101110111011","100110011001","100110011001","101110111011","110011001100","011101110111","011001100110","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011001100110","011101110111","010101010101","010101010101","100110011001","100010001000","011101110111","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011101110111","011101110111","100010001000","100010001000","011001100110","011001100110","100010001000","011101110111","011101110111","011101110111","011001100110","011101110111","010101010101","010101010101","100110011001","100110011001","100010001000","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100010001000","100010001000","100110011001","011101110111","011101110111","011001100110","011001100110","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","010101010101","010101010101","101010101010","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","100110011001","100010001000","100010001000","100110011001","011101110111","011101110111","011001100110","011001100110","011101110111","011101110111","100010001000","100110011001","011101110111","011101110111","010101010101","010101010101","101010101010","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100010001000","100010001000","100110011001","011101110111","100010001000","011001100110","011101110111","010101010101","010101010101","101010101010","101010101010","100010001000","100110011001","011001100110","011001100110","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","100010001000","100010001000","011101110111","100010001000","011001100110","011101110111","010101010101","010101010101","101010101010","101010101010","100010001000","100110011001","011001100110","011001100110","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","100010001000","100010001000","100010001000","011101110111","011101110111","011001100110","011001100110","010101010101","010101010101","101010101010","100110011001","011001100110","011101110111","100010001000","011101110111","011101110111","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100110011001","100110011001","100110011001","100110011001","011101110111","011101110111","011001100110","011001100110","010101010101","010101010101","101010101010","100110011001","011001100110","011001100110","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","010101010101","010101010101","100110011001","100110011001","100010001000","100010001000","100010001000","100110011001","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","100110011001","100110011001","011001100110","011101110111","100010001000","011101110111","011101110111","100010001000","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011101110111","011001100110","011001100110","010101010101","010101010101","100110011001","100110011001","100010001000","100010001000","100010001000","100110011001","011101110111","011101110111","100110011001","100110011001","011101110111","011101110111","100110011001","101010101010","011101110111","011101110111","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011101110111","011101110111","100010001000","100010001000","011001100110","011001100110","100110011001","100110011001","010101010101","011001100110","011101110111","011101110111","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011001100110","011101110111","011101110111","011001100110","011001100110","011101110111","011101110111","100010001000","100110011001","011001100110","011001100110","101110111011","101110111011","011101110111","011001100110","100010001000","100010001000","011101110111","011101110111","011001100110","011001100110","011101110111","011101110111","011001100110","011001100110","011001100110","011001100110","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","011001100110","011001100110","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","011001100110","011001100110","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","010101010101","100010001000");
constant Top: Sprite := ("100010111011","100010111011","100010111010","100010111010","100010111001","100010111001","100111001100","100010111011","100010111011","100010111011","100111001011","100010111011","100010111011","100010111010","011110011001","010001110110","100111001100","101011001100","100111001011","100010111011","011110111010","100010111011","100111001011","100111001011","100010111011","100010111010","100111001011","100111001011","100010111011","101011001100","100111001100","010001110110","100010111011","011010101001","011010101001","011010011000","011010011000","100010111011","100010111011","011110111010","011110101010","011010101001","011110101010","011110101010","011010101001","011010101001","010110000111","010101110111","100111001100","100010111011","100010111011","011110101010","011010101001","011010101001","011010101001","011010101001","010110011000","011010101001","011010101001","011010101001","011010101001","100010111011","011010011001","010001110110","100010111010","011010101001","010110010111","010110010111","100010111011","011110111010","011010111010","011010101001","010110101001","010010010111","010010010111","010110101001","010110101001","010110101001","010010000111","001101100110","100010111011","011010111010","100010111011","011010111010","010110101001","010110011000","010110011000","010110101001","010110101001","010110011000","011010101001","011010101001","011010101001","010110101001","010110011000","010001110110","100010111010","011010101000","010110010111","011110111010","011010111010","011010111010","011010101001","010110101001","010010010111","010010010111","010010010111","010110011000","010110101001","010110011000","011010011001","001101100101","100010111010","011010111010","011010111010","011110111010","011010101001","010110101001","010110011000","010110101001","010110011000","010110010111","011010101001","011010101001","011010111010","011010111001","010110000111","001101100101","100010111010","011010010111","011010101000","011010101000","011010101001","011010101001","010110101001","010010010111","011010101001","010010010111","010010010111","010110011000","100010111010","010110011000","010110001000","010101110111","100010111010","011010101001","011010111010","011010101001","011010101001","010110101001","010110011000","011010101001","011010101001","011010111010","010110010111","010110101000","010110101000","011010101000","010110000111","001101100101","100010111001","011010010111","010110010111","011010101000","010110101001","010110101001","010010010111","011010101001","011110111010","011010101001","010110011000","100010111010","011110111001","011110111010","010110000111","010001110110","100010111010","010110101001","011010101001","011010101001","010110101001","010110101001","010010000111","011010101001","011110111010","011110111010","011010101000","010110010110","010110101000","010110101000","010010000110","001101100101","100010111001","011010010111","010010010111","010010010111","010010010111","010010010111","011010101001","100010111011","011110111010","011010101001","010110010111","011110111001","011110111001","100010111010","011010011000","001101100110","101011001100","010110011000","011010101001","011010101001","011010101001","011010101001","010010000111","011010111010","011110111010","011010101001","010110101000","010110010111","010110010110","010110010111","010001110101","001101100100","100010111001","011010011000","010010010111","010010010111","010010010111","011010101001","011010111010","011110111010","011010111010","010110101001","010010010111","011110111010","100010111010","011110111010","010110011000","010001110110","100010111010","011010101001","011010101001","011010101001","010110011000","010110011000","010110011000","010010000111","011010101001","010110101001","010110010111","010110010111","010110010111","010110010111","010001110110","001101100101","011110101001","011110111010","100010111011","011110111010","010010010111","010010010111","011010101001","011010111010","011010101001","010010010111","010010010111","011010101000","011110111001","011110111001","010110011000","010001110110","100010111010","011010101001","011010101001","010110011000","011110111010","011110111010","011010111010","011010101001","010010011000","010010011000","010110101001","011010111010","011010101001","010110011000","010001110110","001101100100","100111001100","011110111010","011110111010","011010111010","010110011000","010010010111","010110101001","010110101001","010010010111","010110011000","010110011000","010110010111","010110101000","011010101000","010110000111","001101100101","100010111010","011010101001","010110011000","011110111010","100010111011","100010111011","011110111010","011010111010","010110101001","010010011000","011010101001","011110111010","011010111010","010110101001","010010000110","001101100100","100111001100","011110111010","011010111010","011010101001","010110101001","010010010111","010010000111","010010000111","011110111010","011110111010","011110111010","011110111001","010110010111","010110101000","010010000111","001101100101","010010000111","011010101001","011010101001","011110111010","100010111011","011110111010","011010111010","011010101001","010110101001","010110011000","011010101001","011110111010","011010111010","011010101001","010010000111","001101100101","011110011001","011110111010","011010101001","010110101001","010110101001","010010000111","010010010111","011110111010","011110111010","011110111010","011110111010","011110111010","011110111001","010110010111","001101010100","011010011000","010001110110","011010101001","011010111010","100010111011","011110111010","011010111010","011010101001","010110101001","010110101001","010110011000","010110101001","011010111010","011010101001","010110101001","010001100110","001101100101","011110011001","011010001000","011010111010","011010101001","010110101001","010010000111","011110111010","011110111010","011110111010","011110111010","011010101001","011010101001","011010101001","001101100101","100010111011","011110101001","010010000111","001101100110","010110101001","011010111010","011010101001","010110101001","010110101001","010110101001","010010010111","010010010111","010010011000","010110101001","010110101001","010101110111","011110101001","001101100101","011110101010","010001110110","010101110111","011010111010","010010000111","011010101001","011010101001","011110111010","011010101001","011010101001","011010101001","010110101001","001101010101","100010111010","011110101001","011010101001","011010101001","010110011000","010001110110","010110101001","010010010111","010010010111","010010010111","010010010111","011010101001","011110111010","011010101001","010010011000","010101110111","100010111010","010010000111","001101100101","100111001011","011110101010","010110001000","010101110111","011010101001","010110101001","011010101001","011010101001","010110101001","010110101001","010110101001","001101010101","100010111010","011110101010","011010101001","011010111010","011110111010","011110111010","011010011000","010001110110","010110101001","010010010111","011010101001","011110111010","011110111010","011110111010","011010111010","010101110111","100010111010","010110011000","010110001000","010001110110","100111001100","011110111010","011010101001","010110001000","010101110111","010110101001","010110101001","010110101001","010110101001","010010000111","001101010101","100010111010","011110101010","011010111010","011110111010","100010111011","011110111010","011110111010","011110111010","011010011000","001101100110","011110111010","011010111010","011110111010","011110111010","011010111010","010101110111","100010111010","010110011000","011010111010","011110011001","010101110111","100111001011","011110111010","010110101001","010010000111","011010011000","010001110110","010110101001","010010000111","010010000111","001101100110","100010111010","011110101010","011010111010","011110111010","100010111011","011110111010","011110111010","011110111010","011010101001","010110101001","010010000111","010001110110","011010111010","011010111010","011010101001","010101110111","100010111010","010110011000","011010101001","100010111011","011010011001","010101110111","100010111011","011010101001","010110101001","010010000111","011110101001","010110011000","010101110111","010010000111","010001110110","100010111011","011010101001","011010101001","011010101001","011110111010","011110111010","011110111010","011010111010","011010101001","010110101001","010010011000","010110101001","010001110110","001101100110","010110101001","010101110111","100010111010","010110011000","010010000111","011010111010","011110111010","010110011000","010001110110","100010111010","011010101001","011110101001","010010000111","010010000111","011110111010","011010011000","010001110110","100010111011","011010101001","010110101001","010110011000","010110101001","011010101001","011010111010","011010111010","011010101001","010110101001","010010011000","010110011000","010010011000","010110101001","010010000111","001101100110","100010111010","010110011000","010010000111","010010011000","011010101001","011010111010","010110001000","001101100110","100111001100","011110111010","010110011000","011110101001","010010000111","011010101001","011010011000","010001110110","100010111011","011010101001","010010000111","010110011000","010110010111","010110101001","010110101001","010110101001","010010011000","010110011000","010110101001","100010111011","011110111010","011110111010","011010011000","001101100101","100010111010","011010101001","010010011000","010010000111","010010000111","010110101001","010010000111","001101010101","100111001100","011110111010","011010101001","010110101001","010110011000","010110101001","010110000111","010001110110","100010111010","010110011000","010110011000","010110010111","010110010111","010110010111","010110010111","010110010111","010110011000","010110101001","011110111010","011110111010","100010111011","011110111010","010110011000","010001110110","100010111010","011010101001","011110111010","011110111010","010110011000","010110011000","010001110110","001101100101","100111001100","011110111010","011010111010","011010101001","010110011000","010110011000","001101110110","001101010101","011110101001","010110011000","010110010111","011010101000","011110111001","011110111001","010110010111","010110010111","010110011000","010110011000","011010101001","011010111010","011110111010","011010111010","010110001000","010001110110","100010111010","011110111010","100010111011","011110111010","011010111010","010110011000","010001110110","010101110111","100111001011","011110101010","010110101001","010110101001","011110101001","010110011000","010010000111","001101100101","100111001011","100010111010","011010101000","011110111001","011110111001","100010111010","011110111001","011110111001","010110010111","010110011000","010110101001","011010101001","011010101001","011010101001","010010000111","001101100101","100010111010","011110111010","011110111010","100010111011","011110111010","011010101001","010001110110","010001110110","100010111010","011010101001","010110101001","010010000111","010110011000","011010111010","010110011000","010001110110","100111001011","100010111010","010110101000","011010101000","011110111001","011110111001","100010111010","100010111010","011110111001","011010111001","010110011000","010110101001","010110101001","010110101001","010001110110","001101100101","100010111010","100010111011","011110111010","011110111010","011110111010","011010111010","010110001000","001101010101","100111001011","010110011000","010010000111","011110101001","011010111010","011110111010","011110011001","010001110110","100010111011","010110011000","010110101000","010110101000","011110111001","011110111001","011110111001","011110111001","100010111010","100010111010","011010111010","010110011000","010110101001","010110011000","010010000111","001101100110","101011001100","100010111011","011110111010","011110111010","011110111010","011010111010","010010000111","001101100101","011110101001","011110111010","011110101001","011010111010","011110111010","100010111011","011010011000","010001110110","100010111010","010110011000","010110010111","010110101000","010110101000","011010101000","011010101000","011110111001","011010111001","011110111010","100010111011","011110111010","010110011000","010110011000","010010000111","010101110111","101011001100","011110111011","011110111010","011110111010","011010111010","011010101001","010010000111","001101100101","100111001011","011110111010","011010101001","011010111010","011110111010","011010111010","010110011000","010001110110","100010111010","011010101001","010110101001","010110101000","010110010111","010110101000","010110101000","010110101000","011010101001","011010111010","011110111010","011010111010","011010101001","010010000111","010010000111","010101110111","100111001011","011110111011","011110111010","011010111010","011010101001","010110101001","010010000111","001101100101","100111001011","011110111010","011010101001","011110111010","011010111010","011010101001","010110001000","001101100110","100111001011","011110101010","010110101001","010110101001","010110101001","010110010111","010110010111","010110101000","010110101001","010110101001","011010101001","011010111010","011010101001","011010101001","001101110110","001101100101","100010111011","011110111010","011010111010","011010101001","010110101001","010110101001","010001110110","001101100101","100010111010","011110111010","010010000111","011010101001","011010101001","010110101001","010010000111","001101100101","011110111010","011110101010","011010101001","010110101001","010110101001","010110101001","010110101001","010110010111","010110011000","010110011000","010110101001","010110101001","011010101001","010110101001","001101110110","001101100101","100010111010","011110101010","010110101001","010110101001","010110101001","010010011000","001101110110","010001110110","100010111011","011010101001","011110101001","010010000111","010110101001","010110101000","001101110101","001101100101","100111001011","100010111011","011110111010","011010101001","011010101001","010110101001","010110101001","010110101001","010110101001","010110011000","010110011000","010110011000","010110101001","010010011000","001101110110","010001110110","100010111011","011010101001","010110101001","010010011000","010010011000","010010000111","010110011000","010001110110","100010111011","011010011000","010010000111","010001110110","001101110110","010001110110","010001110110","001001010100","100010111010","011010011001","011010011000","010110011000","010110001000","010110001000","010110001000","010110001000","010110001000","010110001000","010001110110","010001110110","010001110110","001101110110","010110011000","010001100110","100010111010","011010011000","010001110110","001101110110","001101110110","010110001000","010110011000","010101110111","011110011001","010001110110","001101100110","001101100101","001101100101","001101100101","001101100101","001101100101","010001110110","010001110110","010001110110","010001110110","010001110110","001101100110","001101100101","001101100101","010001110110","010101110111","010001110110","001101100101","001101010101","010001110110","010101110111","010101110111","010001110110","010001110110","001001010100","001001010100","001101100101","010001110110","010101110111","010101110111");
constant SkyObs : Sprite := ("100101010100","100101010011","100101010100","101001010100","100101010100","100101010100","100001010011","101010011001","100101010100","101001010100","100001000011","101001010100","100101010100","101001010100","100101010100","100101010100","100101010100","100101010011","100101010100","101001010100","100101010100","100101010100","100001010011","101010011001","100101010100","101001010100","100001000011","101001010100","100101010100","101001010100","100101010100","100101010100","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101110101001","101001010100","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","100001000011","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","010100110010","101110101001","101001010100","100001000011","011101000011","011101000011","100001000011","100001000011","100001000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","100001000011","011101000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","101010011001","101001010100","100001000011","011101000011","100001000011","100001000011","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","010100110010","100001000011","100001000011","010100110010","010100110010","010100110010","010100110010","101110011001","101001010100","010100110010","010100110010","011101000011","010100110010","100001000011","010100110010","011101000011","011101000011","010100110010","011101000011","011101000011","011101000011","010100110010","010100110010","101110101001","101001010100","010100110010","010100110010","010100110010","100001000011","010100110010","100001000011","010100110010","101010001000","101010001000","100110001000","100110001000","100110001000","100110001000","101110011001","101110011001","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101010001000","101010001000","100110001000","100110001000","101110101001","101110101001","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101010011000","101010011000","100101010100","101001010100","100001000011","101001010100","100101010100","101001010100","100101010100","100101010100","101001010100","100101010100","100101010011","100101010100","101001010100","100101010100","100101010100","101010011001","101001010100","100101010100","101001010100","100001000011","101001010100","100101010100","101001010100","100101010100","100101010100","100101010100","100101010011","100101010100","101001010100","100101010100","100101010100","101010011001","101001010100","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","100001000011","011101000011","100001000011","100001000011","100001000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","010100110010","101110011001","101001010100","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","011101000011","011101000011","100001000011","011101000011","100001000011","011101000011","011101000011","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","101110011001","101001010100","100001000011","011101000011","100001000011","100001000011","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","101110101001","101001010100","011101000011","100001000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101110101001","101001010100","011101000011","100001000011","011101000011","011101000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","010100110010","101010011001","101001010100","011101000011","100001000011","010100110010","010100110010","100001000011","100001000011","010100110010","011101000011","011101000011","010100110010","010100110010","011101000011","010100110010","010100110010","101110011001","101001010100","010100110010","010100110010","011101000011","010100110010","100001000011","010100110010","011101000011","011101000011","010100110010","011101000011","011101000011","010100110010","011101000011","010100110010","101110011001","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101010001000","101010001000","100110001000","100110001000","101110011001","101110011001","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101110011001","101110011001","100101010100","100101010011","100101010100","101001010100","100101010100","100101010100","100001010011","101010011001","100101010100","101001010100","100001000011","100101010100","100101010011","100101010100","100101010100","100101010100","100101010100","100001010011","101001010100","100101010100","101001010100","100001000011","100001010011","101010011001","101001010100","100101010100","100101010100","101001010100","100101010100","101001010100","100101010100","100101010100","011101000011","100001000011","011101000011","011101000011","100001000011","100001000011","011101000011","101010011001","101001010100","011101000011","011101000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","100001000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","010100110010","101010011001","101001010100","100001000011","011101000011","100001000011","011101000011","100001000011","011101000011","011101000011","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","100001000011","011101000011","011101000011","101110101001","101001010100","011101000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","100001000011","101010011001","101001010100","011101000011","100001000011","100001000011","011101000011","011101000011","100001000011","011101000011","011101000011","100001000011","011101000011","100001000011","011101000011","011101000011","010100110010","101110101001","101001010100","011101000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","010100110010","010100110010","010100110010","010100110010","010100110010","010100110010","010100110010","101110011001","101001010100","011101000011","100001000011","011101000011","010100110010","011101000011","011101000011","010100110010","011101000011","011101000011","010100110010","011101000011","011101000011","010100110010","010100110010","101110101001","101001010100","010100110010","010100110010","010100110010","010100110010","010100110010","010100110010","010100110010","100110001000","100110001000","100110001000","100110001000","100110000111","100110000111","101110011001","101110011001","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101110101001","101110101001","100110001000","100110001000","101010001000","101010001000","100110001000","100110001000","100110001000","100110001000","100101010100","100101010011","100101010100","101001010100","100101010100","100101010100","100001010011","101001010100","100101010100","101001010100","100001000011","101001010100","100101010100","101001010100","100101010100","101010011001","100101010100","100101010011","100101010100","100101010100","100001010011","101001010100","100101010100","101001010100","100001000011","101001010100","100101010100","101001010100","100101010100","100101010100","100101010100","101110101001","101001010100","100001000011","011101000011","011101000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","100001000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101110101001","101001010100","100001000011","011101000011","100001000011","100001000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","100001000011","011101000011","011101000011","011101000011","011101000011","100001000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","100001000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","101010011001","101001010100","011101000011","011101000011","100001000011","100001000011","011101000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","101110011001","101001010100","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","100001000011","100001000011","100001000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","100001000011","011101000011","011101000011","011101000011","010100110010","101110011001","101001010100","011101000011","100001000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","011101000011","010100110010","101010011001","101001010100","010100110010","010100110010","011101000011","011101000011","011101000011","010100110010","011101000011","011101000011","011101000011","010100110010","010100110010","010100110010","010100110010","010100110010","101110011001","101001010100","010100110010","010100110010","100001000011","100001000011","010100110010","011101000011","011101000011","011101000011","010100110010","011101000011","011101000011","010100110010","010100110010","010100110010","101010011001","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101110011001","101110011001","101010001000","101010001000","100110001000","100110001000","100110001000","100110001000","100110001000","100110001000","101010001000","101010001000","100110001000","100110001000","100110001000","100110001000","101010011001","101010011001");
constant FloorObs : Sprite := ("101001010000","101001010000","110101110001","110101110001","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","111010010001","111010010001","111010010001","111010010001","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111010010001","110101110001","110101110001","111010010001","111010010001","111010010001","111010010001","111010010001","111010010001","111010010001","110101110001","101001010000","110101110001","110101110001","111010010001","111010010001","111111010011","111111010011","111010010001","111010010001","110101110001","110101110001","101001010000","110101110001","111010010001","110101110001","110101110001","101001010000","101001010000","111010100100","111010100100","111010010001","111010010001","111010010001","111010010001","111010010001","111111110011","111111110011","111010010001","111111010011","111111010011","111010010001","111010010001","101001010000","110101110001","111010010001","111010010001","111111010011","111111010011","111111010011","111111010011","111010010001","111010010001","111010010001","101001010000","110101110001","111010010001","111010010001","110101110001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111010010001","111111010011","111010110001","111010110001","111111110011","111111110011","111111110011","111111010011","111111010011","111010010001","111010010001","111010010001","111010010001","111111010011","111111111001","111111111001","111111110011","111111110011","111111010011","111111010011","111010010001","111010010001","110101110001","110101110001","111010010001","110101110001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111111010011","111010110001","111010110001","001000000000","001000000000","001000000000","001000000000","111111111001","111111111001","111111010011","111010010001","111010010001","111111010011","111111111001","111111111001","001000000000","001000000000","111010110001","111010110001","111111010011","111111010011","111010010001","101001010000","110101110001","111010010001","110101110001","101001010000","101001010000","101001010000","110101110001","111010010001","111010010001","111111010011","111010110001","001000000000","001000000000","001000000000","001000000000","001000000000","001000000000","111111111001","111111111001","111111010011","111010010001","111111111001","111111111001","001000000000","001000000000","001000000000","001000000000","111010110001","111010110001","111111010011","111111010011","111010010001","111010010001","111010010001","111010010001","101001010000","101001010000","101001010000","110101110001","111010010001","111111010011","111010110001","111010110001","001000000000","001000000000","101010100011","101110100011","101110100011","001000000000","001000000000","111111111001","111111010011","111010010001","111111111001","001000000000","001000000000","101110110011","101110110011","001000000000","001000000000","111010110001","111010110001","111111010011","111111010011","111010010001","111010010001","111010010001","101001010000","101001010000","101001010000","110101110001","111010010001","111111010011","111010110001","111010110001","001000000000","001000000000","101110100011","101110100011","101110100011","101110100011","001000000000","111111111001","111010010001","111010010001","111010110001","001000000000","001000000000","101110110011","101110110011","101110110011","001000000000","001000000000","111111110011","111111110011","111111010011","111111010011","111010010001","111010010001","101001010000","101001010000","101001010000","110101110001","111010010001","111111010011","111010110001","001000000000","001000000000","101110100011","101110100011","101110100011","101110100011","101110110011","101110110011","111010110001","111010010001","111010010001","111010110001","001000000000","001000000000","101110110011","101110110011","101110110011","101110110011","001000000000","001000000000","111111110011","111111110011","111111010011","111010010001","111010010001","101001010000","101001010000","101001010000","110101110001","111010010001","111111010011","111010110001","001000000000","001000000000","101110100011","101110100011","101110100011","101110110011","101110110011","101110110011","111010110001","111010010001","111010010001","111010110001","001000000000","001000000000","101110110011","101110110011","101110110011","101110110011","101110110011","001000000000","001000000000","111111110011","111111010011","111111010011","111010010001","101001010000","101001010000","101001010000","110101110001","111010010001","111010010001","111111110011","001000000000","001000000000","101110110011","101110110011","101110110011","101110110011","101110110011","101110110011","111010110001","111010010001","111010010001","111010110001","001000000000","001000000000","110011000011","110011000011","101110110011","101110110011","101110110011","101110110011","001000000000","001000000000","111010110001","111111010011","111010010001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111111110011","001000000000","001000000000","101110110011","101110110011","101110110011","101110110011","101110110011","110011000011","111010110001","111010010001","111010010001","111010110001","001000000000","001000000000","110011000011","110011000011","110011000011","110011000011","101110110011","101110110011","101110110011","001000000000","111010110001","111111010011","111010010001","101001010000","101001010000","101001010000","111010100100","111010100100","111010010001","111010110001","001000000000","001000000000","101110110011","101110110011","101110110011","110011000011","110011000011","110011000011","111010110001","111010010001","111010010001","111010110001","001000000000","001000000000","110011000011","110011000011","110011000011","110011000011","110011000011","101111000011","101110110011","101110110011","111010110001","111111010011","111010010001","101001010000","101001010000","101001010000","111010100100","111010100100","111010010001","111010110001","001000000000","001000000000","101110110011","101111000011","110011000011","110011000011","110011000011","110011000011","111111110011","111010010001","111010010001","111010110001","001000000000","001000000000","110011000011","110011000011","110011000011","110011000011","110011000011","110011000011","110011000011","101110110011","111010110001","111111010011","111010010001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111010110001","111010110001","001000000000","110011000011","110011000011","110011000011","110011000011","110011000011","111111110011","111111110011","111010010001","111010010001","111010110001","111010110001","001000000000","001000000000","110011000011","110011000011","110011000011","110011000011","110011000011","110011000011","110011000011","111010110001","111111010011","111010010001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111010010001","111010110001","111010110001","001000000000","110011000011","110011000011","110011000011","111111110011","111111110011","111010010001","111010010001","111010010001","111010010001","111010110001","111010110001","001000000000","110011010011","110011000011","110011000011","110011000011","110011000011","110011000011","111111110011","111010110001","111010010001","111010010001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111010010001","111010010001","111010110001","111010110001","111010110001","111010110001","111111110011","111111110011","111010010001","111010010001","111010010001","111010010001","111010010001","111010010001","111010110001","111010110001","111010110001","111010110001","111010110001","111111110011","111010110001","111010110001","111111110011","111010010001","111010010001","110101110001","101001010000","101001010000","101001010000","111010100100","111010010001","111010010001","111111010011","111010110001","111111110011","111111110011","111010010001","111010110001","111010110001","111010110001","111010010001","111010010001","111111110011","111111110011","111010110001","111010010001","111010010001","111010010001","111010110001","111010110001","111010110001","111010010001","111010010001","111010110001","111010110001","111010110001","111010010001","110101110001","101001010000","101001010000","101001010000","111010010001","111010010001","111111010011","111010110001","111010110001","001000000000","111111110011","111111110011","111010110001","001000000000","111010110001","111010110001","111111110011","111111110011","001000000000","111010110001","111010110001","111010010001","111010110001","111010110001","001000000000","111010110001","111010110001","111010110001","111111110011","001000000000","111010110001","111010110001","110101110001","101001010000","101001010000","101001010000","111010010001","111111010011","111010110001","111010110001","001000000000","001000000000","001000000000","111010110001","001000000000","001000000000","001000000000","111010110001","111111110011","001000000000","001000000000","001000000000","111010110001","111010110001","111010110001","001000000000","001000000000","001000000000","111111110011","111111110011","001000000000","001000000000","001000000000","111010110001","110101110001","101001010000","101001010000","101001010000","111010010001","111111110011","111111110011","001000000000","001000000000","110011000011","001000000000","001000000000","001000000000","110011010100","001000000000","001000000000","001000000000","001000000000","110111110100","001000000000","001000000000","001000000000","001000000000","001000000000","110011010100","001000000000","001000000000","001000000000","001000000000","101110110011","001000000000","111010110001","101001010000","101001010000","101001010000","101001010000","111010010001","111111110011","001000000000","001000000000","101111000011","110011000011","110011000011","001000000000","110011010100","110011010100","110111100100","001000000000","001000000000","110111100100","110111100100","110111100100","001000000000","001000000000","001000000000","110111100100","110011010100","110011010100","001000000000","001000000000","110011000011","101110110011","101110110011","001000000000","111010110001","101001010000","101001010000","110101110001","111010010001","111111110011","001000000000","001000000000","101110110011","101111000011","110011000011","110011000011","110011010100","110011010100","110111010100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110111010100","110011010100","110011010100","110011000011","110011000011","110011000011","101110110011","101110110011","101110110011","111010110001","101001010000","101001010000","110101110001","111010010001","111010110001","111010110001","001000000000","001000000000","101110110011","110011000011","110011000011","110011010011","110011010100","110011010100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110011010100","110011010100","110011010011","110011000011","110011000011","110011000011","101110110011","101110110011","101110110011","111111010011","101001010000","101001010000","110101110001","111010010001","111010010001","111010110001","111010110001","001000000000","101110110011","101111000011","110011000011","110011000011","110011010100","110011010100","110011010100","110111100100","110111100100","110111100100","110111100100","110111100100","110111100100","110011010100","110011010100","110011010100","110011010011","110011000011","110011000011","101110110011","101110110011","101110110011","101110110011","111111010011","101001010000","101001010000","110101110001","101001010000","111010010001","111010010001","111010110001","001000000000","101110110011","101110110011","110011000011","111111010011","110011010011","110011010100","110011010100","110011010100","110111100100","111111010011","111010010001","110111100100","110011010100","110011010100","110011010100","110011010011","110011000011","111111010011","110011000011","101110110011","101110110011","101110110011","101110110011","111010110001","101001010000","101001010000","110101110001","101001010000","110101110001","111010010001","111010110001","001000000000","101110110011","101110110011","111111010011","111010010001","110011000011","110011010100","110011010100","110011010100","111010110001","111010010001","111010010001","111010110001","110011010100","110011010100","110011010100","110011010011","110011000011","111111010011","111010010001","101110110011","101110110011","101110110011","111111010011","101001010000","101001010000","101001010000","110101110001","101001010000","110101110001","111010010001","111010110001","001000000000","001000000000","111010110001","111111010011","111010010001","111111010011","110011010011","110011010100","111111010011","110101110001","111010100100","111010010001","111010010001","111010010001","111111010011","111111010011","110011000011","110011000011","111010110001","111010010001","110101110001","101001010000","111010010001","110101110001","101001010000","101001010000","101001010000","101001010000","110101110001","110101110001","111010010001","111010010001","111010110001","111010010001","110101110001","101001010000","111010010001","111010010001","111111010011","111010110001","101001010000","110101110001","111010100100","111010100100","111010010001","110101110001","110101110001","101001010000","111010110001","111010110001","111010010001","111010010001","111010010001","101001010000","111010010001","110101110001","110101110001","101001010000","101001010000","101001010000","110101110001","111010010001","111010010001","111010010001","111010010001","110101110001","110101110001","101001010000","110101110001","111010010001","111010010001","110101110001","110101110001","101001010000","111010100100","111010100100","110101110001","110101110001","101001010000","110101110001","110101110001","111010010001","111010010001","111010010001","110101110001","101001010000","111010010001","111010010001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","111010010001","111010010001","110101110001","110101110001","110101110001","101001010000","110101110001","110101110001","111010010001","110101110001","110101110001","101001010000","110101110001","111010100100","110101110001","101001010000","110101110001","110101110001","111010010001","111010010001","111010010001","110101110001","110101110001","101001010000","110101110001","110101110001","110101110001","101001010000","101001010000","101001010000","110101110001","110101110001","110101110001","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","110101110001","110101110001","101001010000","101001010000","110101110001","110101110001","110101110001","101001010000");
constant Player : Sprite := ("011111000110","011111000110","011111000110","011111000110","011111000110","011010110101","011010110101","011111010110","011111000110","100011000110","011111000110","100011010111","100011000111","100011000111","011111000110","011111000110","100011000111","100011000110","011111000110","011010110101","011010110101","011010110101","011111000101","011111000110","011111000110","011111000110","100011000110","100011000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011010110101","011010110101","011010110100","011010110100","011111000110","011111000110","011011000110","011111000110","100011000111","011111000110","011111000110","011111000110","100011000111","100011000111","011010110101","011010110101","011010110101","011010110101","011010100101","011011000101","011111000110","011111000110","100011010111","100011000110","011111000110","100011000111","011111000110","100011000110","011111000110","011111000110","100011010110","011111010110","011010110101","011010110101","011010110101","011010110101","011111010110","011111000110","011111000110","011111000110","011111010110","011111000110","011111010110","011111000110","011111000110","100011010110","011010110101","011010110100","011010110101","011010110101","011010110101","011010110101","011111010110","011111000110","100011010111","100011000111","100011000111","100011000111","100011000111","011111000110","011111000110","011111000110","011111010110","100011010111","011111010110","011010110101","011010110101","011111000110","100011010110","011111000110","011111000110","011111000110","011111000110","011111010110","011111000110","011111000110","100011000110","100011000110","011111000110","011010110101","011010110101","011010110101","011010110101","011111000110","011111000110","100011000110","100011010111","100011010111","100011000110","100011000110","011111000110","100011000111","100011000111","011111000110","100011010110","011111010110","011111000110","011111000110","100011000110","100011000110","011111010110","011111000110","011010110101","011010110101","011011000101","011111000110","100011000110","100011000110","011011000101","011111000110","011111000110","011111000110","011111010110","011111010110","011111000110","100011000111","100011000111","100011000111","100011000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","100011000111","011111010110","100011000111","011111000110","100011000111","100011000110","100011010111","011110110110","011110110101","011010110101","011010110101","011010110100","011010110101","100011010111","011111000101","011111000110","011011000101","011111010110","011111000110","100011010110","011111000110","011111000110","011111000110","011111010110","100011000111","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","100011000110","100011000111","100011010111","011111010110","100011010111","100011010111","011010110101","011010110101","011010110101","011011000101","011010110101","011111000110","011111000110","011111000101","011111000110","011111010110","100011010110","011111010110","011111010110","100011010110","011111010110","011111000110","011111010110","011111000110","011010110101","011010110101","011111000110","100011010110","100011010110","011111000110","011111000110","011111000110","100011000110","100011010111","100011010111","011111010110","011111000110","100011010111","100011010111","011010110101","011010110101","011010110101","011111000110","011111000110","011111000110","011111000110","011111010110","100011010110","011111010110","011111010110","011111010110","011111000110","011111000110","011111010110","011111000110","011010110101","011010110101","011010110101","011010110101","100011010110","100011000110","100011010110","011111000110","011111000110","011111000110","011111000110","011111010110","100011010110","100011000110","011111000110","011111000110","011111000110","011111000110","011111010110","100011010110","011111000110","011111000110","011111000110","100011010110","100011000110","100011010110","011111000110","011111000110","011111000110","100011000110","011111000110","100011010111","011010110101","011010110101","011010110101","010110110100","011111000110","011111000110","011111000110","100011010111","100011000110","011111000110","011111000110","011111000101","100011010110","100011000110","011111000110","011111000110","011111000110","011111000110","011111010110","100011010110","011111010110","100011000111","011111000110","011111000110","100011010111","011111000110","011111000110","100011000110","011111000110","100011010111","011111010110","100011010111","011111000110","011010110101","011010110101","011111010110","100011010110","100011010110","100011000111","100011010111","011111010110","011111000110","011111000110","011111000110","100011010110","011111000110","100011000110","011111000110","011111000110","011111000110","011111000110","011111010110","011111010110","100011010110","011111000110","011111000110","011111000110","011111000110","011111000110","011010110101","011111000101","011111000110","011111000110","011111000110","011111000110","011111010110","011111000110","011111000110","100011010110","100011010110","100011010111","100011000111","011111000110","011111010110","100011010110","011111000110","100011000110","100011000110","011111000110","100011010110","011111000110","011111000110","011111000110","011111000110","100011010110","011111000110","011111000110","011111000110","011111000110","011111000110","011010110101","011010110101","011010110101","011110110101","011111010110","100011010110","011111000110","011111010110","100011000110","100011010110","011111010110","011111010110","100011000111","100011010110","011111000110","011111000110","011111010110","011010110101","011010110100","100011000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011110110110","011111000110","100011000111","011111000110","011111000110","011010110100","011010110100","011010110101","011010110101","100011010110","100011010110","011111000110","011111000110","100011000110","011111000110","011111000110","100011010110","011111000110","011111000110","011111010110","011111010110","011010110100","011010110100","011010110101","011010110100","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","100011010110","011111000110","100011000110","100011000110","011111000110","011111000110","011111000110","011010110100","011010110101","100011010110","100011000110","100011000110","100011010110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111010110","011111010110","011111000110","011010110101","011010110100","011010110101","011011000101","011111000110","011111000110","011111000110","011111000110","100011000110","100011000110","100011000110","011011000101","011010110100","011111000110","011111000110","011111000110","011111000110","100011000111","100011010111","100011010111","100011010110","100011010110","011111000110","100011010110","011111010101","011111010110","011111010110","011111010110","011111010110","011111010110","011111000110","011111000110","011111000101","011010110101","011010110101","011111000110","011111000110","011111000110","011111000110","011111000110","100011010111","100011010110","011010110101","011010110101","011010110101","011010110100","011111000110","011111000110","100011000111","100011000111","100011010111","100011010110","100011000110","100011010110","100011010110","100011010110","011111010110","011111010110","011111010110","011111000110","100011010111","100011000111","011111000110","011111000110","011111000110","011111000101","100011010111","100011010111","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011010110101","011010110101","011010110101","011010110101","011111000110","100011000110","100011010110","011111000110","011111000110","011111000110","011111000110","100011010110","011111000110","011111000110","011111010110","011010110101","011010110101","011111010110","100011010111","100011010110","100011010110","011111000110","011111000110","011111000110","100011010110","100011000111","011111000110","011111000110","011111000110","011111010110","011111000110","011111000110","100011000110","011010110101","011010100100","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","011010110101","011010110101","011010110101","011010110100","100011010111","100011010111","100011010110","011111000110","011111000110","011111000110","100011000111","011111000110","011111000110","011111000111","011111000110","011111000110","011111010110","100011010111","011111000110","011111000110","011110110110","011110110110","011111000110","011111000110","100011000110","011111000110","011111000110","011111000110","011111000110","100011010111","100011010111","100011000110","011010110101","011010110101","011010110101","011010110101","100011010111","100011010111","100011000110","100011010110","011111000110","100011000111","100011000111","100011000111","011111000110","100011000111","011111000110","100011010110","100011010111","100011010111","100011010111","100011010111","011111000110","011111000110","100011000111","100011000110","100011000110","100011000110","011111000110","011111000110","100011010111","100011010111","100011000111","100011010111","011010110101","011010110101","011010110101","011010110101","100011010111","100011010111","011010110101","100011010111","100011000110","011111000110","100011000111","100011000110","011111000110","011111000110","100011010111","011111000110","011111010110","011111000110","100011000111","100011000110","011111000110","100011000110","100011010110","100011010111","100011010110","100011010111","011111000110","011111000110","100011010110","011111010110","011111010110","011111010110","011010110101","011010110101","011010110101","011010110101","100011010111","011010110101","011010110101","011010110101","011111000110","011111000110","100011010111","011111000110","011111000110","011111000110","011111000110","100011010111","011111010110","011111000110","011111000110","100011000110","011111000110","011111000110","100011010111","100011010111","100011000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111010110","011111010110","011111010110","011010110101","011011000101","011111010110","011110110101","011110110101","011010110101","011010110100","100011010111","100011010110","011111000110","100011000110","011111000110","011111000110","100011000110","100011010110","100011010110","011111000110","100011010110","100011010110","100011010110","011011000101","011010110101","100011010110","011111010110","011111000110","011111010110","100011010110","011111010110","011111010110","100011010110","100011000110","011111010110","011111000110","011111000110","011111000110","100011010110","011110110101","011010110101","011010110101","011010110101","100011010111","100011000110","100011000110","100011010110","011111000110","100011010110","100011000110","100011010110","100011010110","100011010110","011111000110","011011000101","011010110101","011110110101","011010110101","011111010110","011111000110","011111010110","011111000110","011111010110","100011010110","011111000110","100011000110","100011000110","011111010110","011111000110","011111010110","011110110110","011111000110","100011010111","011010110101","100011010111","011111000110","100011010111","011111000110","011111000110","011010110100","011110110101","100011010110","011111000110","100011010111","011111000110","011111010110","011010110101","011010110101","011010110101","011010110101","100011000111","100011000110","011111000110","011010110101","011010110101","100011000110","100011010110","011111000110","011111000110","100011000110","011111000110","011111010110","011110110110","011111000110","011111000110","100011000111","011111000110","100011000111","011111000110","011111000110","011010110101","011010110101","011010110101","011010110101","100011010111","100011010110","011111010110","100011010110","100011010110","011010110101","011010110101","011111000110","100011000110","100011000110","011010110101","011010110101","011111000101","011010110101","011111000110","011111000110","100011000111","011111000110","011111010110","011111000110","011111000110","011111000110","100011010110","011111000110","011111000110","011111000110","011111000110","011111000110","011011000101","011011000101","011010110101","011010110101","011111010110","011111010110","011111000110","100011000111","100011010110","011111010110","011111000110","011111000110","100011000110","011111000110","011010110101","011010110101","011010110101","011010110101","100011010110","100011000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","100011010110","011111000110","011111000110","100011000110","100011000110","011111010110","011111000101","011011000101","011010110101","011010110101","011111010110","011111010110","100011000111","100011000111","100011010111","011111000110","011111000110","011111000110","011111010110","011111010110","011111000110","011010110101","011010110101","100011000110","011111000110","011111000110","011111000110","011111000110","011111000110","011111000110","100011010111","100011010110","011111000110","011111000110","011111000110","100011010111","011111000110","011111000110","100011010110","011010110100","011010110101","011010110101","100011010110","100011010111","011111000110","100011000111","100011000111","100011000111","011111000110","100011010111","100011010110","011111000110","011111000110","011111000110","100011010110","100011010110","011111000110","011111000110","011111000110","011010100101","011010110101","011111000110","100011010111","100011010110","011111000110","011111000110","100011010111","100011010111","100011000110","011111000110","100011010110","100011010110","011110110101","100011010110","100011010111","100011010111","011111010110","011111000110","100011000111","100011010111","100011010111","100011010111","100011010111","011111000110","011111000110","011111000110","011111010110","011111000110","100011000110","011111000110","011010110101","011010110101","011010110101","011010110101","100011000110","011111000110","100011010111","100011010111","100011000111","011111000110","011111000110","011111000110","011111010110","011111000110","100011010110","011111000110","011111000110","100011010111","100011000110","011111000110","100011000111","100011000110","100011010111","100011000110","011111010110","011111010110","011111000110","011111000110","011111000110","100011000110","100011010111","011111000110","011010110101","011010110101","011010110101","011010110101","011111000110","011111000110","100011010111","100011010110","100011010111","100011000111","011111000110","011111000110","011111000110","011111010110","011111000110","011111000110","011111010110","100011010111","100011010111","100011000110","100011000110","100011000110","100011000111","100011000110","100011000110","011111000110","011111000110","100011000110","100011000110","100011000110","100011000110","011111000110","011111000110","011010110101","011010110101","011111000110");



end package ROMS;

package body ROMS is

end package body ROMS;